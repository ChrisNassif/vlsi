module tensor_core_register_file (
	clock_in,
	non_bulk_write_enable_in,
	non_bulk_write_register_address_in,
	non_bulk_write_data_in,
	bulk_write_enable_in,
	bulk_write_data_in,
	read_data_out
);
	reg _sv2v_0;
	parameter NUMBER_OF_REGISTERS = 32;
	input wire clock_in;
	input wire non_bulk_write_enable_in;
	input wire [$clog2(NUMBER_OF_REGISTERS) - 1:0] non_bulk_write_register_address_in;
	input wire [7:0] non_bulk_write_data_in;
	input wire bulk_write_enable_in;
	input wire [(((0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? ((1 - (((NUMBER_OF_REGISTERS - 1) / 16) + 0)) * 4) + (((((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4) - 1) : ((((NUMBER_OF_REGISTERS - 1) / 16) + 1) * 4) - 1) >= (0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? (((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4 : 0) ? ((((0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? ((1 - (((NUMBER_OF_REGISTERS - 1) / 16) + 0)) * 4) + (((((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4) - 1) : ((((NUMBER_OF_REGISTERS - 1) / 16) + 1) * 4) - 1) - (0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? (((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4 : 0)) + 1) * 4) + (((0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? (((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4 : 0) * 4) - 1) : ((((0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? (((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4 : 0) - (0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? ((1 - (((NUMBER_OF_REGISTERS - 1) / 16) + 0)) * 4) + (((((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4) - 1) : ((((NUMBER_OF_REGISTERS - 1) / 16) + 1) * 4) - 1)) + 1) * 4) + (((0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? ((1 - (((NUMBER_OF_REGISTERS - 1) / 16) + 0)) * 4) + (((((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4) - 1) : ((((NUMBER_OF_REGISTERS - 1) / 16) + 1) * 4) - 1) * 4) - 1)) >= ((0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? ((1 - (((NUMBER_OF_REGISTERS - 1) / 16) + 0)) * 4) + (((((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4) - 1) : ((((NUMBER_OF_REGISTERS - 1) / 16) + 1) * 4) - 1) >= (0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? (((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4 : 0) ? (0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? (((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4 : 0) * 4 : (0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? ((1 - (((NUMBER_OF_REGISTERS - 1) / 16) + 0)) * 4) + (((((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4) - 1) : ((((NUMBER_OF_REGISTERS - 1) / 16) + 1) * 4) - 1) * 4) ? (((((0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? ((1 - (((NUMBER_OF_REGISTERS - 1) / 16) + 0)) * 4) + (((((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4) - 1) : ((((NUMBER_OF_REGISTERS - 1) / 16) + 1) * 4) - 1) >= (0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? (((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4 : 0) ? ((((0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? ((1 - (((NUMBER_OF_REGISTERS - 1) / 16) + 0)) * 4) + (((((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4) - 1) : ((((NUMBER_OF_REGISTERS - 1) / 16) + 1) * 4) - 1) - (0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? (((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4 : 0)) + 1) * 4) + (((0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? (((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4 : 0) * 4) - 1) : ((((0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? (((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4 : 0) - (0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? ((1 - (((NUMBER_OF_REGISTERS - 1) / 16) + 0)) * 4) + (((((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4) - 1) : ((((NUMBER_OF_REGISTERS - 1) / 16) + 1) * 4) - 1)) + 1) * 4) + (((0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? ((1 - (((NUMBER_OF_REGISTERS - 1) / 16) + 0)) * 4) + (((((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4) - 1) : ((((NUMBER_OF_REGISTERS - 1) / 16) + 1) * 4) - 1) * 4) - 1)) - ((0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? ((1 - (((NUMBER_OF_REGISTERS - 1) / 16) + 0)) * 4) + (((((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4) - 1) : ((((NUMBER_OF_REGISTERS - 1) / 16) + 1) * 4) - 1) >= (0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? (((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4 : 0) ? (0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? (((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4 : 0) * 4 : (0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? ((1 - (((NUMBER_OF_REGISTERS - 1) / 16) + 0)) * 4) + (((((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4) - 1) : ((((NUMBER_OF_REGISTERS - 1) / 16) + 1) * 4) - 1) * 4)) + 1) * 8) + ((((0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? ((1 - (((NUMBER_OF_REGISTERS - 1) / 16) + 0)) * 4) + (((((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4) - 1) : ((((NUMBER_OF_REGISTERS - 1) / 16) + 1) * 4) - 1) >= (0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? (((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4 : 0) ? (0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? (((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4 : 0) * 4 : (0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? ((1 - (((NUMBER_OF_REGISTERS - 1) / 16) + 0)) * 4) + (((((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4) - 1) : ((((NUMBER_OF_REGISTERS - 1) / 16) + 1) * 4) - 1) * 4) * 8) - 1) : (((((0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? ((1 - (((NUMBER_OF_REGISTERS - 1) / 16) + 0)) * 4) + (((((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4) - 1) : ((((NUMBER_OF_REGISTERS - 1) / 16) + 1) * 4) - 1) >= (0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? (((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4 : 0) ? (0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? (((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4 : 0) * 4 : (0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? ((1 - (((NUMBER_OF_REGISTERS - 1) / 16) + 0)) * 4) + (((((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4) - 1) : ((((NUMBER_OF_REGISTERS - 1) / 16) + 1) * 4) - 1) * 4) - ((0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? ((1 - (((NUMBER_OF_REGISTERS - 1) / 16) + 0)) * 4) + (((((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4) - 1) : ((((NUMBER_OF_REGISTERS - 1) / 16) + 1) * 4) - 1) >= (0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? (((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4 : 0) ? ((((0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? ((1 - (((NUMBER_OF_REGISTERS - 1) / 16) + 0)) * 4) + (((((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4) - 1) : ((((NUMBER_OF_REGISTERS - 1) / 16) + 1) * 4) - 1) - (0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? (((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4 : 0)) + 1) * 4) + (((0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? (((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4 : 0) * 4) - 1) : ((((0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? (((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4 : 0) - (0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? ((1 - (((NUMBER_OF_REGISTERS - 1) / 16) + 0)) * 4) + (((((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4) - 1) : ((((NUMBER_OF_REGISTERS - 1) / 16) + 1) * 4) - 1)) + 1) * 4) + (((0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? ((1 - (((NUMBER_OF_REGISTERS - 1) / 16) + 0)) * 4) + (((((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4) - 1) : ((((NUMBER_OF_REGISTERS - 1) / 16) + 1) * 4) - 1) * 4) - 1))) + 1) * 8) + ((((0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? ((1 - (((NUMBER_OF_REGISTERS - 1) / 16) + 0)) * 4) + (((((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4) - 1) : ((((NUMBER_OF_REGISTERS - 1) / 16) + 1) * 4) - 1) >= (0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? (((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4 : 0) ? ((((0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? ((1 - (((NUMBER_OF_REGISTERS - 1) / 16) + 0)) * 4) + (((((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4) - 1) : ((((NUMBER_OF_REGISTERS - 1) / 16) + 1) * 4) - 1) - (0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? (((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4 : 0)) + 1) * 4) + (((0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? (((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4 : 0) * 4) - 1) : ((((0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? (((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4 : 0) - (0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? ((1 - (((NUMBER_OF_REGISTERS - 1) / 16) + 0)) * 4) + (((((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4) - 1) : ((((NUMBER_OF_REGISTERS - 1) / 16) + 1) * 4) - 1)) + 1) * 4) + (((0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? ((1 - (((NUMBER_OF_REGISTERS - 1) / 16) + 0)) * 4) + (((((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4) - 1) : ((((NUMBER_OF_REGISTERS - 1) / 16) + 1) * 4) - 1) * 4) - 1)) * 8) - 1)):(((0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? ((1 - (((NUMBER_OF_REGISTERS - 1) / 16) + 0)) * 4) + (((((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4) - 1) : ((((NUMBER_OF_REGISTERS - 1) / 16) + 1) * 4) - 1) >= (0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? (((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4 : 0) ? ((((0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? ((1 - (((NUMBER_OF_REGISTERS - 1) / 16) + 0)) * 4) + (((((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4) - 1) : ((((NUMBER_OF_REGISTERS - 1) / 16) + 1) * 4) - 1) - (0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? (((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4 : 0)) + 1) * 4) + (((0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? (((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4 : 0) * 4) - 1) : ((((0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? (((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4 : 0) - (0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? ((1 - (((NUMBER_OF_REGISTERS - 1) / 16) + 0)) * 4) + (((((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4) - 1) : ((((NUMBER_OF_REGISTERS - 1) / 16) + 1) * 4) - 1)) + 1) * 4) + (((0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? ((1 - (((NUMBER_OF_REGISTERS - 1) / 16) + 0)) * 4) + (((((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4) - 1) : ((((NUMBER_OF_REGISTERS - 1) / 16) + 1) * 4) - 1) * 4) - 1)) >= ((0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? ((1 - (((NUMBER_OF_REGISTERS - 1) / 16) + 0)) * 4) + (((((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4) - 1) : ((((NUMBER_OF_REGISTERS - 1) / 16) + 1) * 4) - 1) >= (0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? (((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4 : 0) ? (0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? (((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4 : 0) * 4 : (0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? ((1 - (((NUMBER_OF_REGISTERS - 1) / 16) + 0)) * 4) + (((((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4) - 1) : ((((NUMBER_OF_REGISTERS - 1) / 16) + 1) * 4) - 1) * 4) ? ((0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? ((1 - (((NUMBER_OF_REGISTERS - 1) / 16) + 0)) * 4) + (((((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4) - 1) : ((((NUMBER_OF_REGISTERS - 1) / 16) + 1) * 4) - 1) >= (0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? (((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4 : 0) ? (0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? (((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4 : 0) * 4 : (0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? ((1 - (((NUMBER_OF_REGISTERS - 1) / 16) + 0)) * 4) + (((((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4) - 1) : ((((NUMBER_OF_REGISTERS - 1) / 16) + 1) * 4) - 1) * 4) * 8 : ((0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? ((1 - (((NUMBER_OF_REGISTERS - 1) / 16) + 0)) * 4) + (((((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4) - 1) : ((((NUMBER_OF_REGISTERS - 1) / 16) + 1) * 4) - 1) >= (0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? (((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4 : 0) ? ((((0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? ((1 - (((NUMBER_OF_REGISTERS - 1) / 16) + 0)) * 4) + (((((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4) - 1) : ((((NUMBER_OF_REGISTERS - 1) / 16) + 1) * 4) - 1) - (0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? (((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4 : 0)) + 1) * 4) + (((0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? (((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4 : 0) * 4) - 1) : ((((0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? (((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4 : 0) - (0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? ((1 - (((NUMBER_OF_REGISTERS - 1) / 16) + 0)) * 4) + (((((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4) - 1) : ((((NUMBER_OF_REGISTERS - 1) / 16) + 1) * 4) - 1)) + 1) * 4) + (((0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? ((1 - (((NUMBER_OF_REGISTERS - 1) / 16) + 0)) * 4) + (((((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4) - 1) : ((((NUMBER_OF_REGISTERS - 1) / 16) + 1) * 4) - 1) * 4) - 1)) * 8)] bulk_write_data_in;
	output reg [(((0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? ((1 - (((NUMBER_OF_REGISTERS - 1) / 16) + 0)) * 4) + (((((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4) - 1) : ((((NUMBER_OF_REGISTERS - 1) / 16) + 1) * 4) - 1) >= (0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? (((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4 : 0) ? ((((0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? ((1 - (((NUMBER_OF_REGISTERS - 1) / 16) + 0)) * 4) + (((((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4) - 1) : ((((NUMBER_OF_REGISTERS - 1) / 16) + 1) * 4) - 1) - (0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? (((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4 : 0)) + 1) * 4) + (((0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? (((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4 : 0) * 4) - 1) : ((((0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? (((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4 : 0) - (0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? ((1 - (((NUMBER_OF_REGISTERS - 1) / 16) + 0)) * 4) + (((((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4) - 1) : ((((NUMBER_OF_REGISTERS - 1) / 16) + 1) * 4) - 1)) + 1) * 4) + (((0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? ((1 - (((NUMBER_OF_REGISTERS - 1) / 16) + 0)) * 4) + (((((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4) - 1) : ((((NUMBER_OF_REGISTERS - 1) / 16) + 1) * 4) - 1) * 4) - 1)) >= ((0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? ((1 - (((NUMBER_OF_REGISTERS - 1) / 16) + 0)) * 4) + (((((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4) - 1) : ((((NUMBER_OF_REGISTERS - 1) / 16) + 1) * 4) - 1) >= (0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? (((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4 : 0) ? (0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? (((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4 : 0) * 4 : (0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? ((1 - (((NUMBER_OF_REGISTERS - 1) / 16) + 0)) * 4) + (((((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4) - 1) : ((((NUMBER_OF_REGISTERS - 1) / 16) + 1) * 4) - 1) * 4) ? (((((0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? ((1 - (((NUMBER_OF_REGISTERS - 1) / 16) + 0)) * 4) + (((((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4) - 1) : ((((NUMBER_OF_REGISTERS - 1) / 16) + 1) * 4) - 1) >= (0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? (((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4 : 0) ? ((((0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? ((1 - (((NUMBER_OF_REGISTERS - 1) / 16) + 0)) * 4) + (((((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4) - 1) : ((((NUMBER_OF_REGISTERS - 1) / 16) + 1) * 4) - 1) - (0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? (((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4 : 0)) + 1) * 4) + (((0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? (((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4 : 0) * 4) - 1) : ((((0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? (((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4 : 0) - (0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? ((1 - (((NUMBER_OF_REGISTERS - 1) / 16) + 0)) * 4) + (((((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4) - 1) : ((((NUMBER_OF_REGISTERS - 1) / 16) + 1) * 4) - 1)) + 1) * 4) + (((0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? ((1 - (((NUMBER_OF_REGISTERS - 1) / 16) + 0)) * 4) + (((((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4) - 1) : ((((NUMBER_OF_REGISTERS - 1) / 16) + 1) * 4) - 1) * 4) - 1)) - ((0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? ((1 - (((NUMBER_OF_REGISTERS - 1) / 16) + 0)) * 4) + (((((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4) - 1) : ((((NUMBER_OF_REGISTERS - 1) / 16) + 1) * 4) - 1) >= (0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? (((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4 : 0) ? (0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? (((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4 : 0) * 4 : (0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? ((1 - (((NUMBER_OF_REGISTERS - 1) / 16) + 0)) * 4) + (((((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4) - 1) : ((((NUMBER_OF_REGISTERS - 1) / 16) + 1) * 4) - 1) * 4)) + 1) * 8) + ((((0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? ((1 - (((NUMBER_OF_REGISTERS - 1) / 16) + 0)) * 4) + (((((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4) - 1) : ((((NUMBER_OF_REGISTERS - 1) / 16) + 1) * 4) - 1) >= (0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? (((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4 : 0) ? (0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? (((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4 : 0) * 4 : (0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? ((1 - (((NUMBER_OF_REGISTERS - 1) / 16) + 0)) * 4) + (((((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4) - 1) : ((((NUMBER_OF_REGISTERS - 1) / 16) + 1) * 4) - 1) * 4) * 8) - 1) : (((((0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? ((1 - (((NUMBER_OF_REGISTERS - 1) / 16) + 0)) * 4) + (((((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4) - 1) : ((((NUMBER_OF_REGISTERS - 1) / 16) + 1) * 4) - 1) >= (0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? (((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4 : 0) ? (0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? (((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4 : 0) * 4 : (0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? ((1 - (((NUMBER_OF_REGISTERS - 1) / 16) + 0)) * 4) + (((((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4) - 1) : ((((NUMBER_OF_REGISTERS - 1) / 16) + 1) * 4) - 1) * 4) - ((0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? ((1 - (((NUMBER_OF_REGISTERS - 1) / 16) + 0)) * 4) + (((((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4) - 1) : ((((NUMBER_OF_REGISTERS - 1) / 16) + 1) * 4) - 1) >= (0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? (((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4 : 0) ? ((((0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? ((1 - (((NUMBER_OF_REGISTERS - 1) / 16) + 0)) * 4) + (((((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4) - 1) : ((((NUMBER_OF_REGISTERS - 1) / 16) + 1) * 4) - 1) - (0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? (((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4 : 0)) + 1) * 4) + (((0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? (((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4 : 0) * 4) - 1) : ((((0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? (((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4 : 0) - (0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? ((1 - (((NUMBER_OF_REGISTERS - 1) / 16) + 0)) * 4) + (((((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4) - 1) : ((((NUMBER_OF_REGISTERS - 1) / 16) + 1) * 4) - 1)) + 1) * 4) + (((0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? ((1 - (((NUMBER_OF_REGISTERS - 1) / 16) + 0)) * 4) + (((((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4) - 1) : ((((NUMBER_OF_REGISTERS - 1) / 16) + 1) * 4) - 1) * 4) - 1))) + 1) * 8) + ((((0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? ((1 - (((NUMBER_OF_REGISTERS - 1) / 16) + 0)) * 4) + (((((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4) - 1) : ((((NUMBER_OF_REGISTERS - 1) / 16) + 1) * 4) - 1) >= (0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? (((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4 : 0) ? ((((0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? ((1 - (((NUMBER_OF_REGISTERS - 1) / 16) + 0)) * 4) + (((((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4) - 1) : ((((NUMBER_OF_REGISTERS - 1) / 16) + 1) * 4) - 1) - (0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? (((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4 : 0)) + 1) * 4) + (((0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? (((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4 : 0) * 4) - 1) : ((((0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? (((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4 : 0) - (0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? ((1 - (((NUMBER_OF_REGISTERS - 1) / 16) + 0)) * 4) + (((((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4) - 1) : ((((NUMBER_OF_REGISTERS - 1) / 16) + 1) * 4) - 1)) + 1) * 4) + (((0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? ((1 - (((NUMBER_OF_REGISTERS - 1) / 16) + 0)) * 4) + (((((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4) - 1) : ((((NUMBER_OF_REGISTERS - 1) / 16) + 1) * 4) - 1) * 4) - 1)) * 8) - 1)):(((0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? ((1 - (((NUMBER_OF_REGISTERS - 1) / 16) + 0)) * 4) + (((((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4) - 1) : ((((NUMBER_OF_REGISTERS - 1) / 16) + 1) * 4) - 1) >= (0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? (((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4 : 0) ? ((((0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? ((1 - (((NUMBER_OF_REGISTERS - 1) / 16) + 0)) * 4) + (((((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4) - 1) : ((((NUMBER_OF_REGISTERS - 1) / 16) + 1) * 4) - 1) - (0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? (((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4 : 0)) + 1) * 4) + (((0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? (((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4 : 0) * 4) - 1) : ((((0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? (((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4 : 0) - (0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? ((1 - (((NUMBER_OF_REGISTERS - 1) / 16) + 0)) * 4) + (((((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4) - 1) : ((((NUMBER_OF_REGISTERS - 1) / 16) + 1) * 4) - 1)) + 1) * 4) + (((0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? ((1 - (((NUMBER_OF_REGISTERS - 1) / 16) + 0)) * 4) + (((((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4) - 1) : ((((NUMBER_OF_REGISTERS - 1) / 16) + 1) * 4) - 1) * 4) - 1)) >= ((0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? ((1 - (((NUMBER_OF_REGISTERS - 1) / 16) + 0)) * 4) + (((((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4) - 1) : ((((NUMBER_OF_REGISTERS - 1) / 16) + 1) * 4) - 1) >= (0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? (((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4 : 0) ? (0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? (((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4 : 0) * 4 : (0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? ((1 - (((NUMBER_OF_REGISTERS - 1) / 16) + 0)) * 4) + (((((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4) - 1) : ((((NUMBER_OF_REGISTERS - 1) / 16) + 1) * 4) - 1) * 4) ? ((0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? ((1 - (((NUMBER_OF_REGISTERS - 1) / 16) + 0)) * 4) + (((((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4) - 1) : ((((NUMBER_OF_REGISTERS - 1) / 16) + 1) * 4) - 1) >= (0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? (((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4 : 0) ? (0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? (((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4 : 0) * 4 : (0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? ((1 - (((NUMBER_OF_REGISTERS - 1) / 16) + 0)) * 4) + (((((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4) - 1) : ((((NUMBER_OF_REGISTERS - 1) / 16) + 1) * 4) - 1) * 4) * 8 : ((0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? ((1 - (((NUMBER_OF_REGISTERS - 1) / 16) + 0)) * 4) + (((((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4) - 1) : ((((NUMBER_OF_REGISTERS - 1) / 16) + 1) * 4) - 1) >= (0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? (((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4 : 0) ? ((((0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? ((1 - (((NUMBER_OF_REGISTERS - 1) / 16) + 0)) * 4) + (((((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4) - 1) : ((((NUMBER_OF_REGISTERS - 1) / 16) + 1) * 4) - 1) - (0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? (((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4 : 0)) + 1) * 4) + (((0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? (((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4 : 0) * 4) - 1) : ((((0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? (((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4 : 0) - (0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? ((1 - (((NUMBER_OF_REGISTERS - 1) / 16) + 0)) * 4) + (((((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4) - 1) : ((((NUMBER_OF_REGISTERS - 1) / 16) + 1) * 4) - 1)) + 1) * 4) + (((0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? ((1 - (((NUMBER_OF_REGISTERS - 1) / 16) + 0)) * 4) + (((((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4) - 1) : ((((NUMBER_OF_REGISTERS - 1) / 16) + 1) * 4) - 1) * 4) - 1)) * 8)] read_data_out;
	reg [7:0] registers [0:((NUMBER_OF_REGISTERS - 1) / 16) + 0][0:3][0:3];
	always @(*) begin
		if (_sv2v_0)
			;
		begin : sv2v_autoblock_1
			reg signed [31:0] n;
			for (n = 0; n < 2; n = n + 1)
				begin : sv2v_autoblock_2
					reg signed [31:0] i;
					for (i = 0; i < 4; i = i + 1)
						begin : sv2v_autoblock_3
							reg signed [31:0] j;
							for (j = 0; j < 4; j = j + 1)
								read_data_out[(((0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? ((1 - (((NUMBER_OF_REGISTERS - 1) / 16) + 0)) * 4) + (((((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4) - 1) : ((((NUMBER_OF_REGISTERS - 1) / 16) + 1) * 4) - 1) >= (0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? (((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4 : 0) ? ((((0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? ((1 - (((NUMBER_OF_REGISTERS - 1) / 16) + 0)) * 4) + (((((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4) - 1) : ((((NUMBER_OF_REGISTERS - 1) / 16) + 1) * 4) - 1) - (0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? (((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4 : 0)) + 1) * 4) + (((0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? (((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4 : 0) * 4) - 1) : ((((0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? (((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4 : 0) - (0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? ((1 - (((NUMBER_OF_REGISTERS - 1) / 16) + 0)) * 4) + (((((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4) - 1) : ((((NUMBER_OF_REGISTERS - 1) / 16) + 1) * 4) - 1)) + 1) * 4) + (((0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? ((1 - (((NUMBER_OF_REGISTERS - 1) / 16) + 0)) * 4) + (((((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4) - 1) : ((((NUMBER_OF_REGISTERS - 1) / 16) + 1) * 4) - 1) * 4) - 1)) >= ((0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? ((1 - (((NUMBER_OF_REGISTERS - 1) / 16) + 0)) * 4) + (((((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4) - 1) : ((((NUMBER_OF_REGISTERS - 1) / 16) + 1) * 4) - 1) >= (0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? (((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4 : 0) ? (0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? (((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4 : 0) * 4 : (0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? ((1 - (((NUMBER_OF_REGISTERS - 1) / 16) + 0)) * 4) + (((((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4) - 1) : ((((NUMBER_OF_REGISTERS - 1) / 16) + 1) * 4) - 1) * 4) ? (((0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? ((1 - (((NUMBER_OF_REGISTERS - 1) / 16) + 0)) * 4) + (((((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4) - 1) : ((((NUMBER_OF_REGISTERS - 1) / 16) + 1) * 4) - 1) >= (0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? (((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4 : 0) ? ((0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? n : (((NUMBER_OF_REGISTERS - 1) / 16) + 0) - n) * 4) + (3 - i) : (0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? (((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4 : 0) - ((((0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? n : (((NUMBER_OF_REGISTERS - 1) / 16) + 0) - n) * 4) + (3 - i)) - (0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? ((1 - (((NUMBER_OF_REGISTERS - 1) / 16) + 0)) * 4) + (((((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4) - 1) : ((((NUMBER_OF_REGISTERS - 1) / 16) + 1) * 4) - 1))) * 4) + (3 - j) : ((0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? ((1 - (((NUMBER_OF_REGISTERS - 1) / 16) + 0)) * 4) + (((((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4) - 1) : ((((NUMBER_OF_REGISTERS - 1) / 16) + 1) * 4) - 1) >= (0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? (((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4 : 0) ? (0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? (((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4 : 0) * 4 : (0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? ((1 - (((NUMBER_OF_REGISTERS - 1) / 16) + 0)) * 4) + (((((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4) - 1) : ((((NUMBER_OF_REGISTERS - 1) / 16) + 1) * 4) - 1) * 4) - (((((0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? ((1 - (((NUMBER_OF_REGISTERS - 1) / 16) + 0)) * 4) + (((((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4) - 1) : ((((NUMBER_OF_REGISTERS - 1) / 16) + 1) * 4) - 1) >= (0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? (((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4 : 0) ? ((0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? n : (((NUMBER_OF_REGISTERS - 1) / 16) + 0) - n) * 4) + (3 - i) : (0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? (((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4 : 0) - ((((0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? n : (((NUMBER_OF_REGISTERS - 1) / 16) + 0) - n) * 4) + (3 - i)) - (0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? ((1 - (((NUMBER_OF_REGISTERS - 1) / 16) + 0)) * 4) + (((((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4) - 1) : ((((NUMBER_OF_REGISTERS - 1) / 16) + 1) * 4) - 1))) * 4) + (3 - j)) - ((0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? ((1 - (((NUMBER_OF_REGISTERS - 1) / 16) + 0)) * 4) + (((((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4) - 1) : ((((NUMBER_OF_REGISTERS - 1) / 16) + 1) * 4) - 1) >= (0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? (((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4 : 0) ? ((((0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? ((1 - (((NUMBER_OF_REGISTERS - 1) / 16) + 0)) * 4) + (((((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4) - 1) : ((((NUMBER_OF_REGISTERS - 1) / 16) + 1) * 4) - 1) - (0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? (((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4 : 0)) + 1) * 4) + (((0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? (((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4 : 0) * 4) - 1) : ((((0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? (((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4 : 0) - (0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? ((1 - (((NUMBER_OF_REGISTERS - 1) / 16) + 0)) * 4) + (((((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4) - 1) : ((((NUMBER_OF_REGISTERS - 1) / 16) + 1) * 4) - 1)) + 1) * 4) + (((0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? ((1 - (((NUMBER_OF_REGISTERS - 1) / 16) + 0)) * 4) + (((((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4) - 1) : ((((NUMBER_OF_REGISTERS - 1) / 16) + 1) * 4) - 1) * 4) - 1)))) * 8+:8] = registers[n][i][j];
						end
				end
		end
	end
	initial begin : sv2v_autoblock_4
		reg signed [31:0] i;
		for (i = 0; i < (((NUMBER_OF_REGISTERS - 1) / 16) + 1); i = i + 1)
			begin : sv2v_autoblock_5
				reg signed [31:0] j;
				for (j = 0; j < 4; j = j + 1)
					begin : sv2v_autoblock_6
						reg signed [31:0] k;
						for (k = 0; k < 4; k = k + 1)
							registers[i][j][k] = 8'b00000000;
					end
			end
	end
	always @(posedge clock_in)
		if (bulk_write_enable_in) begin : sv2v_autoblock_7
			reg signed [31:0] i;
			for (i = 0; i < (((NUMBER_OF_REGISTERS - 1) / 16) + 1); i = i + 1)
				begin : sv2v_autoblock_8
					reg signed [31:0] j;
					for (j = 0; j < 4; j = j + 1)
						begin : sv2v_autoblock_9
							reg signed [31:0] k;
							for (k = 0; k < 4; k = k + 1)
								registers[i][j][k] <= bulk_write_data_in[(((0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? ((1 - (((NUMBER_OF_REGISTERS - 1) / 16) + 0)) * 4) + (((((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4) - 1) : ((((NUMBER_OF_REGISTERS - 1) / 16) + 1) * 4) - 1) >= (0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? (((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4 : 0) ? ((((0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? ((1 - (((NUMBER_OF_REGISTERS - 1) / 16) + 0)) * 4) + (((((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4) - 1) : ((((NUMBER_OF_REGISTERS - 1) / 16) + 1) * 4) - 1) - (0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? (((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4 : 0)) + 1) * 4) + (((0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? (((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4 : 0) * 4) - 1) : ((((0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? (((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4 : 0) - (0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? ((1 - (((NUMBER_OF_REGISTERS - 1) / 16) + 0)) * 4) + (((((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4) - 1) : ((((NUMBER_OF_REGISTERS - 1) / 16) + 1) * 4) - 1)) + 1) * 4) + (((0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? ((1 - (((NUMBER_OF_REGISTERS - 1) / 16) + 0)) * 4) + (((((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4) - 1) : ((((NUMBER_OF_REGISTERS - 1) / 16) + 1) * 4) - 1) * 4) - 1)) >= ((0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? ((1 - (((NUMBER_OF_REGISTERS - 1) / 16) + 0)) * 4) + (((((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4) - 1) : ((((NUMBER_OF_REGISTERS - 1) / 16) + 1) * 4) - 1) >= (0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? (((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4 : 0) ? (0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? (((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4 : 0) * 4 : (0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? ((1 - (((NUMBER_OF_REGISTERS - 1) / 16) + 0)) * 4) + (((((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4) - 1) : ((((NUMBER_OF_REGISTERS - 1) / 16) + 1) * 4) - 1) * 4) ? (((0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? ((1 - (((NUMBER_OF_REGISTERS - 1) / 16) + 0)) * 4) + (((((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4) - 1) : ((((NUMBER_OF_REGISTERS - 1) / 16) + 1) * 4) - 1) >= (0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? (((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4 : 0) ? ((0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? i : (((NUMBER_OF_REGISTERS - 1) / 16) + 0) - i) * 4) + (3 - j) : (0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? (((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4 : 0) - ((((0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? i : (((NUMBER_OF_REGISTERS - 1) / 16) + 0) - i) * 4) + (3 - j)) - (0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? ((1 - (((NUMBER_OF_REGISTERS - 1) / 16) + 0)) * 4) + (((((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4) - 1) : ((((NUMBER_OF_REGISTERS - 1) / 16) + 1) * 4) - 1))) * 4) + (3 - k) : ((0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? ((1 - (((NUMBER_OF_REGISTERS - 1) / 16) + 0)) * 4) + (((((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4) - 1) : ((((NUMBER_OF_REGISTERS - 1) / 16) + 1) * 4) - 1) >= (0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? (((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4 : 0) ? (0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? (((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4 : 0) * 4 : (0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? ((1 - (((NUMBER_OF_REGISTERS - 1) / 16) + 0)) * 4) + (((((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4) - 1) : ((((NUMBER_OF_REGISTERS - 1) / 16) + 1) * 4) - 1) * 4) - (((((0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? ((1 - (((NUMBER_OF_REGISTERS - 1) / 16) + 0)) * 4) + (((((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4) - 1) : ((((NUMBER_OF_REGISTERS - 1) / 16) + 1) * 4) - 1) >= (0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? (((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4 : 0) ? ((0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? i : (((NUMBER_OF_REGISTERS - 1) / 16) + 0) - i) * 4) + (3 - j) : (0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? (((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4 : 0) - ((((0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? i : (((NUMBER_OF_REGISTERS - 1) / 16) + 0) - i) * 4) + (3 - j)) - (0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? ((1 - (((NUMBER_OF_REGISTERS - 1) / 16) + 0)) * 4) + (((((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4) - 1) : ((((NUMBER_OF_REGISTERS - 1) / 16) + 1) * 4) - 1))) * 4) + (3 - k)) - ((0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? ((1 - (((NUMBER_OF_REGISTERS - 1) / 16) + 0)) * 4) + (((((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4) - 1) : ((((NUMBER_OF_REGISTERS - 1) / 16) + 1) * 4) - 1) >= (0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? (((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4 : 0) ? ((((0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? ((1 - (((NUMBER_OF_REGISTERS - 1) / 16) + 0)) * 4) + (((((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4) - 1) : ((((NUMBER_OF_REGISTERS - 1) / 16) + 1) * 4) - 1) - (0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? (((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4 : 0)) + 1) * 4) + (((0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? (((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4 : 0) * 4) - 1) : ((((0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? (((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4 : 0) - (0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? ((1 - (((NUMBER_OF_REGISTERS - 1) / 16) + 0)) * 4) + (((((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4) - 1) : ((((NUMBER_OF_REGISTERS - 1) / 16) + 1) * 4) - 1)) + 1) * 4) + (((0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? ((1 - (((NUMBER_OF_REGISTERS - 1) / 16) + 0)) * 4) + (((((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4) - 1) : ((((NUMBER_OF_REGISTERS - 1) / 16) + 1) * 4) - 1) * 4) - 1)))) * 8+:8];
						end
				end
		end
		else if (non_bulk_write_enable_in)
			registers[non_bulk_write_register_address_in / 16][(non_bulk_write_register_address_in % 16) / 4][non_bulk_write_register_address_in % 4] <= non_bulk_write_data_in;
	genvar _gv_i_1;
	genvar _gv_j_1;
	genvar _gv_k_1;
	generate
		for (_gv_i_1 = 0; _gv_i_1 < (((NUMBER_OF_REGISTERS - 1) / 16) + 1); _gv_i_1 = _gv_i_1 + 1) begin : expose_regs1
			localparam i = _gv_i_1;
			for (_gv_j_1 = 0; _gv_j_1 < 4; _gv_j_1 = _gv_j_1 + 1) begin : expose_regs2
				localparam j = _gv_j_1;
				for (_gv_k_1 = 0; _gv_k_1 < 4; _gv_k_1 = _gv_k_1 + 1) begin : expose_regs3
					localparam k = _gv_k_1;
					wire [7:0] reg_wire = registers[i][j][k];
					wire [7:0] read_data_out_ = read_data_out[(((0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? ((1 - (((NUMBER_OF_REGISTERS - 1) / 16) + 0)) * 4) + (((((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4) - 1) : ((((NUMBER_OF_REGISTERS - 1) / 16) + 1) * 4) - 1) >= (0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? (((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4 : 0) ? ((((0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? ((1 - (((NUMBER_OF_REGISTERS - 1) / 16) + 0)) * 4) + (((((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4) - 1) : ((((NUMBER_OF_REGISTERS - 1) / 16) + 1) * 4) - 1) - (0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? (((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4 : 0)) + 1) * 4) + (((0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? (((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4 : 0) * 4) - 1) : ((((0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? (((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4 : 0) - (0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? ((1 - (((NUMBER_OF_REGISTERS - 1) / 16) + 0)) * 4) + (((((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4) - 1) : ((((NUMBER_OF_REGISTERS - 1) / 16) + 1) * 4) - 1)) + 1) * 4) + (((0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? ((1 - (((NUMBER_OF_REGISTERS - 1) / 16) + 0)) * 4) + (((((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4) - 1) : ((((NUMBER_OF_REGISTERS - 1) / 16) + 1) * 4) - 1) * 4) - 1)) >= ((0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? ((1 - (((NUMBER_OF_REGISTERS - 1) / 16) + 0)) * 4) + (((((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4) - 1) : ((((NUMBER_OF_REGISTERS - 1) / 16) + 1) * 4) - 1) >= (0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? (((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4 : 0) ? (0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? (((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4 : 0) * 4 : (0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? ((1 - (((NUMBER_OF_REGISTERS - 1) / 16) + 0)) * 4) + (((((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4) - 1) : ((((NUMBER_OF_REGISTERS - 1) / 16) + 1) * 4) - 1) * 4) ? (((0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? ((1 - (((NUMBER_OF_REGISTERS - 1) / 16) + 0)) * 4) + (((((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4) - 1) : ((((NUMBER_OF_REGISTERS - 1) / 16) + 1) * 4) - 1) >= (0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? (((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4 : 0) ? ((0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? i : (((NUMBER_OF_REGISTERS - 1) / 16) + 0) - i) * 4) + (3 - j) : (0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? (((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4 : 0) - ((((0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? i : (((NUMBER_OF_REGISTERS - 1) / 16) + 0) - i) * 4) + (3 - j)) - (0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? ((1 - (((NUMBER_OF_REGISTERS - 1) / 16) + 0)) * 4) + (((((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4) - 1) : ((((NUMBER_OF_REGISTERS - 1) / 16) + 1) * 4) - 1))) * 4) + (3 - k) : ((0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? ((1 - (((NUMBER_OF_REGISTERS - 1) / 16) + 0)) * 4) + (((((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4) - 1) : ((((NUMBER_OF_REGISTERS - 1) / 16) + 1) * 4) - 1) >= (0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? (((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4 : 0) ? (0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? (((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4 : 0) * 4 : (0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? ((1 - (((NUMBER_OF_REGISTERS - 1) / 16) + 0)) * 4) + (((((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4) - 1) : ((((NUMBER_OF_REGISTERS - 1) / 16) + 1) * 4) - 1) * 4) - (((((0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? ((1 - (((NUMBER_OF_REGISTERS - 1) / 16) + 0)) * 4) + (((((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4) - 1) : ((((NUMBER_OF_REGISTERS - 1) / 16) + 1) * 4) - 1) >= (0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? (((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4 : 0) ? ((0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? i : (((NUMBER_OF_REGISTERS - 1) / 16) + 0) - i) * 4) + (3 - j) : (0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? (((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4 : 0) - ((((0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? i : (((NUMBER_OF_REGISTERS - 1) / 16) + 0) - i) * 4) + (3 - j)) - (0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? ((1 - (((NUMBER_OF_REGISTERS - 1) / 16) + 0)) * 4) + (((((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4) - 1) : ((((NUMBER_OF_REGISTERS - 1) / 16) + 1) * 4) - 1))) * 4) + (3 - k)) - ((0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? ((1 - (((NUMBER_OF_REGISTERS - 1) / 16) + 0)) * 4) + (((((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4) - 1) : ((((NUMBER_OF_REGISTERS - 1) / 16) + 1) * 4) - 1) >= (0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? (((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4 : 0) ? ((((0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? ((1 - (((NUMBER_OF_REGISTERS - 1) / 16) + 0)) * 4) + (((((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4) - 1) : ((((NUMBER_OF_REGISTERS - 1) / 16) + 1) * 4) - 1) - (0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? (((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4 : 0)) + 1) * 4) + (((0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? (((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4 : 0) * 4) - 1) : ((((0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? (((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4 : 0) - (0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? ((1 - (((NUMBER_OF_REGISTERS - 1) / 16) + 0)) * 4) + (((((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4) - 1) : ((((NUMBER_OF_REGISTERS - 1) / 16) + 1) * 4) - 1)) + 1) * 4) + (((0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? ((1 - (((NUMBER_OF_REGISTERS - 1) / 16) + 0)) * 4) + (((((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4) - 1) : ((((NUMBER_OF_REGISTERS - 1) / 16) + 1) * 4) - 1) * 4) - 1)))) * 8+:8];
					wire [7:0] bulk_write_data_in_ = bulk_write_data_in[(((0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? ((1 - (((NUMBER_OF_REGISTERS - 1) / 16) + 0)) * 4) + (((((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4) - 1) : ((((NUMBER_OF_REGISTERS - 1) / 16) + 1) * 4) - 1) >= (0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? (((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4 : 0) ? ((((0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? ((1 - (((NUMBER_OF_REGISTERS - 1) / 16) + 0)) * 4) + (((((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4) - 1) : ((((NUMBER_OF_REGISTERS - 1) / 16) + 1) * 4) - 1) - (0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? (((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4 : 0)) + 1) * 4) + (((0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? (((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4 : 0) * 4) - 1) : ((((0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? (((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4 : 0) - (0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? ((1 - (((NUMBER_OF_REGISTERS - 1) / 16) + 0)) * 4) + (((((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4) - 1) : ((((NUMBER_OF_REGISTERS - 1) / 16) + 1) * 4) - 1)) + 1) * 4) + (((0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? ((1 - (((NUMBER_OF_REGISTERS - 1) / 16) + 0)) * 4) + (((((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4) - 1) : ((((NUMBER_OF_REGISTERS - 1) / 16) + 1) * 4) - 1) * 4) - 1)) >= ((0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? ((1 - (((NUMBER_OF_REGISTERS - 1) / 16) + 0)) * 4) + (((((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4) - 1) : ((((NUMBER_OF_REGISTERS - 1) / 16) + 1) * 4) - 1) >= (0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? (((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4 : 0) ? (0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? (((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4 : 0) * 4 : (0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? ((1 - (((NUMBER_OF_REGISTERS - 1) / 16) + 0)) * 4) + (((((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4) - 1) : ((((NUMBER_OF_REGISTERS - 1) / 16) + 1) * 4) - 1) * 4) ? (((0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? ((1 - (((NUMBER_OF_REGISTERS - 1) / 16) + 0)) * 4) + (((((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4) - 1) : ((((NUMBER_OF_REGISTERS - 1) / 16) + 1) * 4) - 1) >= (0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? (((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4 : 0) ? ((0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? i : (((NUMBER_OF_REGISTERS - 1) / 16) + 0) - i) * 4) + (3 - j) : (0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? (((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4 : 0) - ((((0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? i : (((NUMBER_OF_REGISTERS - 1) / 16) + 0) - i) * 4) + (3 - j)) - (0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? ((1 - (((NUMBER_OF_REGISTERS - 1) / 16) + 0)) * 4) + (((((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4) - 1) : ((((NUMBER_OF_REGISTERS - 1) / 16) + 1) * 4) - 1))) * 4) + (3 - k) : ((0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? ((1 - (((NUMBER_OF_REGISTERS - 1) / 16) + 0)) * 4) + (((((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4) - 1) : ((((NUMBER_OF_REGISTERS - 1) / 16) + 1) * 4) - 1) >= (0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? (((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4 : 0) ? (0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? (((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4 : 0) * 4 : (0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? ((1 - (((NUMBER_OF_REGISTERS - 1) / 16) + 0)) * 4) + (((((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4) - 1) : ((((NUMBER_OF_REGISTERS - 1) / 16) + 1) * 4) - 1) * 4) - (((((0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? ((1 - (((NUMBER_OF_REGISTERS - 1) / 16) + 0)) * 4) + (((((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4) - 1) : ((((NUMBER_OF_REGISTERS - 1) / 16) + 1) * 4) - 1) >= (0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? (((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4 : 0) ? ((0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? i : (((NUMBER_OF_REGISTERS - 1) / 16) + 0) - i) * 4) + (3 - j) : (0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? (((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4 : 0) - ((((0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? i : (((NUMBER_OF_REGISTERS - 1) / 16) + 0) - i) * 4) + (3 - j)) - (0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? ((1 - (((NUMBER_OF_REGISTERS - 1) / 16) + 0)) * 4) + (((((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4) - 1) : ((((NUMBER_OF_REGISTERS - 1) / 16) + 1) * 4) - 1))) * 4) + (3 - k)) - ((0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? ((1 - (((NUMBER_OF_REGISTERS - 1) / 16) + 0)) * 4) + (((((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4) - 1) : ((((NUMBER_OF_REGISTERS - 1) / 16) + 1) * 4) - 1) >= (0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? (((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4 : 0) ? ((((0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? ((1 - (((NUMBER_OF_REGISTERS - 1) / 16) + 0)) * 4) + (((((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4) - 1) : ((((NUMBER_OF_REGISTERS - 1) / 16) + 1) * 4) - 1) - (0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? (((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4 : 0)) + 1) * 4) + (((0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? (((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4 : 0) * 4) - 1) : ((((0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? (((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4 : 0) - (0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? ((1 - (((NUMBER_OF_REGISTERS - 1) / 16) + 0)) * 4) + (((((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4) - 1) : ((((NUMBER_OF_REGISTERS - 1) / 16) + 1) * 4) - 1)) + 1) * 4) + (((0 >= (((NUMBER_OF_REGISTERS - 1) / 16) + 0) ? ((1 - (((NUMBER_OF_REGISTERS - 1) / 16) + 0)) * 4) + (((((NUMBER_OF_REGISTERS - 1) / 16) + 0) * 4) - 1) : ((((NUMBER_OF_REGISTERS - 1) / 16) + 1) * 4) - 1) * 4) - 1)))) * 8+:8];
				end
			end
		end
	endgenerate
	initial _sv2v_0 = 0;
endmodule
