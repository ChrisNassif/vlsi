`timescale 1ns / 1ps
`default_nettype wire

module cpu (input logic clock_in, input logic machine_code);


    // always @(posedge clock) begin

    // end

  

endmodule